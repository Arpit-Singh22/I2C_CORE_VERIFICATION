`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "../rtl/i2c_master_top.v"
`include "../common/i2c_if.sv"
//`include "../master/i2c_seq_item.sv"
//`include "../master/i2c_driver.sv"
//`include "../common/i2c_monitor.sv"
//`include "../master/i2c_agent.sv"
`include "../top/i2c_env.sv"
`include "../top/i2c_test.sv"
`include "../top/top.sv"
