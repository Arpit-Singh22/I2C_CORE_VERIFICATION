interface i2c_if (input bit clk, input bit rst_n);
  // Add signals later
endinterface
