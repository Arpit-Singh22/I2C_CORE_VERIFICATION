
`include "uvm_macros.svh"
class i2c_agent extends uvm_agent;
  `uvm_component_utils(i2c_agent)
  i2c_driver drv;
  i2c_monitor mon;
  function new(string name, uvm_component parent); super.new(name, parent); endfunction
  function void build_phase(uvm_phase phase);
    drv = i2c_driver::type_id::create("drv", this);
    mon = i2c_monitor::type_id::create("mon", this);
  endfunction
endclass
