interface i2c_if;
	logic scl;
	tri sda;
endinterface
